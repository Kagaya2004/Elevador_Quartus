// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// Created on Sun Apr 30 14:53:57 2023

// synthesis message_off 10175

`timescale 1ns/1ns

module Mov_Elevador (
    clock,reset,EN,ACT,
    SA0,SA1,SA2);

    input clock;
    input reset;
    input EN;
    input ACT;
    tri0 reset;
    tri0 EN;
    tri0 ACT;
    output SA0;
    output SA1;
    output SA2;
    reg SA0;
    reg SA1;
    reg SA2;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter T=0,A1=1,A2=2,A3=3,A4=4;

    always @(posedge clock or posedge reset)
    begin
        if (reset) begin
            fstate <= T;
        end
        else begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or EN or ACT)
    begin
        SA0 <= 1'b0;
        SA1 <= 1'b0;
        SA2 <= 1'b0;
        case (fstate)
            T: begin
                if ((EN == 1'b0))
                    reg_fstate <= T;
                else if (((ACT == 1'b1) & (EN == 1'b1)))
                    reg_fstate <= A1;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= T;

                SA0 <= 1'b1;

                SA1 <= 1'b0;

                SA2 <= 1'b0;
            end
            A1: begin
                if (((ACT == 1'b0) & (EN == 1'b1)))
                    reg_fstate <= T;
                else if ((EN == 1'b0))
                    reg_fstate <= A1;
                else if (((ACT == 1'b1) & (EN == 1'b1)))
                    reg_fstate <= A2;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= A1;

                SA0 <= 1'b0;

                SA1 <= 1'b1;

                SA2 <= 1'b0;
            end
            A2: begin
                if (((ACT == 1'b0) & (EN == 1'b1)))
                    reg_fstate <= A1;
                else if ((EN == 1'b0))
                    reg_fstate <= A2;
                else if (((ACT == 1'b1) & (EN == 1'b1)))
                    reg_fstate <= A3;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= A2;

                SA0 <= 1'b1;

                SA1 <= 1'b1;

                SA2 <= 1'b0;
            end
            A3: begin
                if (((ACT == 1'b0) & (EN == 1'b1)))
                    reg_fstate <= A2;
                else if ((EN == 1'b0))
                    reg_fstate <= A3;
                else if (((ACT == 1'b1) & (EN == 1'b1)))
                    reg_fstate <= A4;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= A3;

                SA0 <= 1'b0;

                SA1 <= 1'b0;

                SA2 <= 1'b1;
            end
            A4: begin
                if (((ACT == 1'b0) & (EN == 1'b1)))
                    reg_fstate <= A3;
                else if ((EN == 1'b0))
                    reg_fstate <= A4;
                // Inserting 'else' block to prevent latch inference
                else
                    reg_fstate <= A4;

                SA0 <= 1'b1;

                SA1 <= 1'b0;

                SA2 <= 1'b1;
            end
            default: begin
                SA0 <= 1'bx;
                SA1 <= 1'bx;
                SA2 <= 1'bx;
                $display ("Reach undefined state");
            end
        endcase
    end
endmodule // Mov_Elevador
